****************************************************************************************
	
This template defines a block RAM configured in 1024 x 18-bit single port mode and 
conneceted to act as a single port ROM.

****************************************************************************************

The next line is used to determine where the template actually starts and must exist.
{begin template}
--
-- Definition of a single port ROM for KCPSM3 program defined by {name}.psm
--
-- Generated by KCPSM3 Assembler {timestamp}. 
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity {name} is
  Port (
    clk_i           : in  std_logic;
    cke_i           : in  std_logic;
    address_i       : in  std_logic_vector(10-1 downto 0);
    instruction_o   : out std_logic_vector(18-1 downto 0)
    );
end {name};
--
architecture rtl of {name} is

begin

  process (clk_i) is
  begin  -- process
    if rising_edge(clk_i)
    then
      if (cke_i = '1')
      then
        case conv_integer(address_i) is
{CASE_BODY10-instruction_o}
          when others => instruction_o <= (others => '0');
        end case;
      end if;
    end if;
  end process;
  
--
end rtl;


architecture rom of {name} is

  type mem_t is array (0 to 2**10-1) of std_logic_vector(18-1 downto 0);

  signal rom : mem_t :=
    (   0 => "{INITX_000}"
    ,   1 => "{INITX_001}"
    ,   2 => "{INITX_002}"
    ,   3 => "{INITX_003}"
    ,   4 => "{INITX_004}"
    ,   5 => "{INITX_005}"
    ,   6 => "{INITX_006}"
    ,   7 => "{INITX_007}"
    ,   8 => "{INITX_008}"
    ,   9 => "{INITX_009}"
    ,  10 => "{INITX_00a}"
    ,  11 => "{INITX_00b}"
    ,  12 => "{INITX_00c}"
    ,  13 => "{INITX_00d}"
    ,  14 => "{INITX_00e}"
    ,  15 => "{INITX_00f}"
    ,  16 => "{INITX_010}"
    ,  17 => "{INITX_011}"
    ,  18 => "{INITX_012}"
    ,  19 => "{INITX_013}"
    ,  20 => "{INITX_014}"
    ,  21 => "{INITX_015}"
    ,  22 => "{INITX_016}"
    ,  23 => "{INITX_017}"
    ,  24 => "{INITX_018}"
    ,  25 => "{INITX_019}"
    ,  26 => "{INITX_01a}"
    ,  27 => "{INITX_01b}"
    ,  28 => "{INITX_01c}"
    ,  29 => "{INITX_01d}"
    ,  30 => "{INITX_01e}"
    ,  31 => "{INITX_01f}"
    ,  32 => "{INITX_020}"
    ,  33 => "{INITX_021}"
    ,  34 => "{INITX_022}"
    ,  35 => "{INITX_023}"
    ,  36 => "{INITX_024}"
    ,  37 => "{INITX_025}"
    ,  38 => "{INITX_026}"
    ,  39 => "{INITX_027}"
    ,  40 => "{INITX_028}"
    ,  41 => "{INITX_029}"
    ,  42 => "{INITX_02a}"
    ,  43 => "{INITX_02b}"
    ,  44 => "{INITX_02c}"
    ,  45 => "{INITX_02d}"
    ,  46 => "{INITX_02e}"
    ,  47 => "{INITX_02f}"
    ,  48 => "{INITX_030}"
    ,  49 => "{INITX_031}"
    ,  50 => "{INITX_032}"
    ,  51 => "{INITX_033}"
    ,  52 => "{INITX_034}"
    ,  53 => "{INITX_035}"
    ,  54 => "{INITX_036}"
    ,  55 => "{INITX_037}"
    ,  56 => "{INITX_038}"
    ,  57 => "{INITX_039}"
    ,  58 => "{INITX_03a}"
    ,  59 => "{INITX_03b}"
    ,  60 => "{INITX_03c}"
    ,  61 => "{INITX_03d}"
    ,  62 => "{INITX_03e}"
    ,  63 => "{INITX_03f}"
    ,  64 => "{INITX_040}"
    ,  65 => "{INITX_041}"
    ,  66 => "{INITX_042}"
    ,  67 => "{INITX_043}"
    ,  68 => "{INITX_044}"
    ,  69 => "{INITX_045}"
    ,  70 => "{INITX_046}"
    ,  71 => "{INITX_047}"
    ,  72 => "{INITX_048}"
    ,  73 => "{INITX_049}"
    ,  74 => "{INITX_04a}"
    ,  75 => "{INITX_04b}"
    ,  76 => "{INITX_04c}"
    ,  77 => "{INITX_04d}"
    ,  78 => "{INITX_04e}"
    ,  79 => "{INITX_04f}"
    ,  80 => "{INITX_050}"
    ,  81 => "{INITX_051}"
    ,  82 => "{INITX_052}"
    ,  83 => "{INITX_053}"
    ,  84 => "{INITX_054}"
    ,  85 => "{INITX_055}"
    ,  86 => "{INITX_056}"
    ,  87 => "{INITX_057}"
    ,  88 => "{INITX_058}"
    ,  89 => "{INITX_059}"
    ,  90 => "{INITX_05a}"
    ,  91 => "{INITX_05b}"
    ,  92 => "{INITX_05c}"
    ,  93 => "{INITX_05d}"
    ,  94 => "{INITX_05e}"
    ,  95 => "{INITX_05f}"
    ,  96 => "{INITX_060}"
    ,  97 => "{INITX_061}"
    ,  98 => "{INITX_062}"
    ,  99 => "{INITX_063}"
    , 100 => "{INITX_064}"
    , 101 => "{INITX_065}"
    , 102 => "{INITX_066}"
    , 103 => "{INITX_067}"
    , 104 => "{INITX_068}"
    , 105 => "{INITX_069}"
    , 106 => "{INITX_06a}"
    , 107 => "{INITX_06b}"
    , 108 => "{INITX_06c}"
    , 109 => "{INITX_06d}"
    , 110 => "{INITX_06e}"
    , 111 => "{INITX_06f}"
    , 112 => "{INITX_070}"
    , 113 => "{INITX_071}"
    , 114 => "{INITX_072}"
    , 115 => "{INITX_073}"
    , 116 => "{INITX_074}"
    , 117 => "{INITX_075}"
    , 118 => "{INITX_076}"
    , 119 => "{INITX_077}"
    , 120 => "{INITX_078}"
    , 121 => "{INITX_079}"
    , 122 => "{INITX_07a}"
    , 123 => "{INITX_07b}"
    , 124 => "{INITX_07c}"
    , 125 => "{INITX_07d}"
    , 126 => "{INITX_07e}"
    , 127 => "{INITX_07f}"
    , 128 => "{INITX_080}"
    , 129 => "{INITX_081}"
    , 130 => "{INITX_082}"
    , 131 => "{INITX_083}"
    , 132 => "{INITX_084}"
    , 133 => "{INITX_085}"
    , 134 => "{INITX_086}"
    , 135 => "{INITX_087}"
    , 136 => "{INITX_088}"
    , 137 => "{INITX_089}"
    , 138 => "{INITX_08a}"
    , 139 => "{INITX_08b}"
    , 140 => "{INITX_08c}"
    , 141 => "{INITX_08d}"
    , 142 => "{INITX_08e}"
    , 143 => "{INITX_08f}"
    , 144 => "{INITX_090}"
    , 145 => "{INITX_091}"
    , 146 => "{INITX_092}"
    , 147 => "{INITX_093}"
    , 148 => "{INITX_094}"
    , 149 => "{INITX_095}"
    , 150 => "{INITX_096}"
    , 151 => "{INITX_097}"
    , 152 => "{INITX_098}"
    , 153 => "{INITX_099}"
    , 154 => "{INITX_09a}"
    , 155 => "{INITX_09b}"
    , 156 => "{INITX_09c}"
    , 157 => "{INITX_09d}"
    , 158 => "{INITX_09e}"
    , 159 => "{INITX_09f}"
    , 160 => "{INITX_0a0}"
    , 161 => "{INITX_0a1}"
    , 162 => "{INITX_0a2}"
    , 163 => "{INITX_0a3}"
    , 164 => "{INITX_0a4}"
    , 165 => "{INITX_0a5}"
    , 166 => "{INITX_0a6}"
    , 167 => "{INITX_0a7}"
    , 168 => "{INITX_0a8}"
    , 169 => "{INITX_0a9}"
    , 170 => "{INITX_0aa}"
    , 171 => "{INITX_0ab}"
    , 172 => "{INITX_0ac}"
    , 173 => "{INITX_0ad}"
    , 174 => "{INITX_0ae}"
    , 175 => "{INITX_0af}"
    , 176 => "{INITX_0b0}"
    , 177 => "{INITX_0b1}"
    , 178 => "{INITX_0b2}"
    , 179 => "{INITX_0b3}"
    , 180 => "{INITX_0b4}"
    , 181 => "{INITX_0b5}"
    , 182 => "{INITX_0b6}"
    , 183 => "{INITX_0b7}"
    , 184 => "{INITX_0b8}"
    , 185 => "{INITX_0b9}"
    , 186 => "{INITX_0ba}"
    , 187 => "{INITX_0bb}"
    , 188 => "{INITX_0bc}"
    , 189 => "{INITX_0bd}"
    , 190 => "{INITX_0be}"
    , 191 => "{INITX_0bf}"
    , 192 => "{INITX_0c0}"
    , 193 => "{INITX_0c1}"
    , 194 => "{INITX_0c2}"
    , 195 => "{INITX_0c3}"
    , 196 => "{INITX_0c4}"
    , 197 => "{INITX_0c5}"
    , 198 => "{INITX_0c6}"
    , 199 => "{INITX_0c7}"
    , 200 => "{INITX_0c8}"
    , 201 => "{INITX_0c9}"
    , 202 => "{INITX_0ca}"
    , 203 => "{INITX_0cb}"
    , 204 => "{INITX_0cc}"
    , 205 => "{INITX_0cd}"
    , 206 => "{INITX_0ce}"
    , 207 => "{INITX_0cf}"
    , 208 => "{INITX_0d0}"
    , 209 => "{INITX_0d1}"
    , 210 => "{INITX_0d2}"
    , 211 => "{INITX_0d3}"
    , 212 => "{INITX_0d4}"
    , 213 => "{INITX_0d5}"
    , 214 => "{INITX_0d6}"
    , 215 => "{INITX_0d7}"
    , 216 => "{INITX_0d8}"
    , 217 => "{INITX_0d9}"
    , 218 => "{INITX_0da}"
    , 219 => "{INITX_0db}"
    , 220 => "{INITX_0dc}"
    , 221 => "{INITX_0dd}"
    , 222 => "{INITX_0de}"
    , 223 => "{INITX_0df}"
    , 224 => "{INITX_0e0}"
    , 225 => "{INITX_0e1}"
    , 226 => "{INITX_0e2}"
    , 227 => "{INITX_0e3}"
    , 228 => "{INITX_0e4}"
    , 229 => "{INITX_0e5}"
    , 230 => "{INITX_0e6}"
    , 231 => "{INITX_0e7}"
    , 232 => "{INITX_0e8}"
    , 233 => "{INITX_0e9}"
    , 234 => "{INITX_0ea}"
    , 235 => "{INITX_0eb}"
    , 236 => "{INITX_0ec}"
    , 237 => "{INITX_0ed}"
    , 238 => "{INITX_0ee}"
    , 239 => "{INITX_0ef}"
    , 240 => "{INITX_0f0}"
    , 241 => "{INITX_0f1}"
    , 242 => "{INITX_0f2}"
    , 243 => "{INITX_0f3}"
    , 244 => "{INITX_0f4}"
    , 245 => "{INITX_0f5}"
    , 246 => "{INITX_0f6}"
    , 247 => "{INITX_0f7}"
    , 248 => "{INITX_0f8}"
    , 249 => "{INITX_0f9}"
    , 250 => "{INITX_0fa}"
    , 251 => "{INITX_0fb}"
    , 252 => "{INITX_0fc}"
    , 253 => "{INITX_0fd}"
    , 254 => "{INITX_0fe}"
    , 255 => "{INITX_0ff}"
    , 256 => "{INITX_100}"
    , 257 => "{INITX_101}"
    , 258 => "{INITX_102}"
    , 259 => "{INITX_103}"
    , 260 => "{INITX_104}"
    , 261 => "{INITX_105}"
    , 262 => "{INITX_106}"
    , 263 => "{INITX_107}"
    , 264 => "{INITX_108}"
    , 265 => "{INITX_109}"
    , 266 => "{INITX_10a}"
    , 267 => "{INITX_10b}"
    , 268 => "{INITX_10c}"
    , 269 => "{INITX_10d}"
    , 270 => "{INITX_10e}"
    , 271 => "{INITX_10f}"
    , 272 => "{INITX_110}"
    , 273 => "{INITX_111}"
    , 274 => "{INITX_112}"
    , 275 => "{INITX_113}"
    , 276 => "{INITX_114}"
    , 277 => "{INITX_115}"
    , 278 => "{INITX_116}"
    , 279 => "{INITX_117}"
    , 280 => "{INITX_118}"
    , 281 => "{INITX_119}"
    , 282 => "{INITX_11a}"
    , 283 => "{INITX_11b}"
    , 284 => "{INITX_11c}"
    , 285 => "{INITX_11d}"
    , 286 => "{INITX_11e}"
    , 287 => "{INITX_11f}"
    , 288 => "{INITX_120}"
    , 289 => "{INITX_121}"
    , 290 => "{INITX_122}"
    , 291 => "{INITX_123}"
    , 292 => "{INITX_124}"
    , 293 => "{INITX_125}"
    , 294 => "{INITX_126}"
    , 295 => "{INITX_127}"
    , 296 => "{INITX_128}"
    , 297 => "{INITX_129}"
    , 298 => "{INITX_12a}"
    , 299 => "{INITX_12b}"
    , 300 => "{INITX_12c}"
    , 301 => "{INITX_12d}"
    , 302 => "{INITX_12e}"
    , 303 => "{INITX_12f}"
    , 304 => "{INITX_130}"
    , 305 => "{INITX_131}"
    , 306 => "{INITX_132}"
    , 307 => "{INITX_133}"
    , 308 => "{INITX_134}"
    , 309 => "{INITX_135}"
    , 310 => "{INITX_136}"
    , 311 => "{INITX_137}"
    , 312 => "{INITX_138}"
    , 313 => "{INITX_139}"
    , 314 => "{INITX_13a}"
    , 315 => "{INITX_13b}"
    , 316 => "{INITX_13c}"
    , 317 => "{INITX_13d}"
    , 318 => "{INITX_13e}"
    , 319 => "{INITX_13f}"
    , 320 => "{INITX_140}"
    , 321 => "{INITX_141}"
    , 322 => "{INITX_142}"
    , 323 => "{INITX_143}"
    , 324 => "{INITX_144}"
    , 325 => "{INITX_145}"
    , 326 => "{INITX_146}"
    , 327 => "{INITX_147}"
    , 328 => "{INITX_148}"
    , 329 => "{INITX_149}"
    , 330 => "{INITX_14a}"
    , 331 => "{INITX_14b}"
    , 332 => "{INITX_14c}"
    , 333 => "{INITX_14d}"
    , 334 => "{INITX_14e}"
    , 335 => "{INITX_14f}"
    , 336 => "{INITX_150}"
    , 337 => "{INITX_151}"
    , 338 => "{INITX_152}"
    , 339 => "{INITX_153}"
    , 340 => "{INITX_154}"
    , 341 => "{INITX_155}"
    , 342 => "{INITX_156}"
    , 343 => "{INITX_157}"
    , 344 => "{INITX_158}"
    , 345 => "{INITX_159}"
    , 346 => "{INITX_15a}"
    , 347 => "{INITX_15b}"
    , 348 => "{INITX_15c}"
    , 349 => "{INITX_15d}"
    , 350 => "{INITX_15e}"
    , 351 => "{INITX_15f}"
    , 352 => "{INITX_160}"
    , 353 => "{INITX_161}"
    , 354 => "{INITX_162}"
    , 355 => "{INITX_163}"
    , 356 => "{INITX_164}"
    , 357 => "{INITX_165}"
    , 358 => "{INITX_166}"
    , 359 => "{INITX_167}"
    , 360 => "{INITX_168}"
    , 361 => "{INITX_169}"
    , 362 => "{INITX_16a}"
    , 363 => "{INITX_16b}"
    , 364 => "{INITX_16c}"
    , 365 => "{INITX_16d}"
    , 366 => "{INITX_16e}"
    , 367 => "{INITX_16f}"
    , 368 => "{INITX_170}"
    , 369 => "{INITX_171}"
    , 370 => "{INITX_172}"
    , 371 => "{INITX_173}"
    , 372 => "{INITX_174}"
    , 373 => "{INITX_175}"
    , 374 => "{INITX_176}"
    , 375 => "{INITX_177}"
    , 376 => "{INITX_178}"
    , 377 => "{INITX_179}"
    , 378 => "{INITX_17a}"
    , 379 => "{INITX_17b}"
    , 380 => "{INITX_17c}"
    , 381 => "{INITX_17d}"
    , 382 => "{INITX_17e}"
    , 383 => "{INITX_17f}"
    , 384 => "{INITX_180}"
    , 385 => "{INITX_181}"
    , 386 => "{INITX_182}"
    , 387 => "{INITX_183}"
    , 388 => "{INITX_184}"
    , 389 => "{INITX_185}"
    , 390 => "{INITX_186}"
    , 391 => "{INITX_187}"
    , 392 => "{INITX_188}"
    , 393 => "{INITX_189}"
    , 394 => "{INITX_18a}"
    , 395 => "{INITX_18b}"
    , 396 => "{INITX_18c}"
    , 397 => "{INITX_18d}"
    , 398 => "{INITX_18e}"
    , 399 => "{INITX_18f}"
    , 400 => "{INITX_190}"
    , 401 => "{INITX_191}"
    , 402 => "{INITX_192}"
    , 403 => "{INITX_193}"
    , 404 => "{INITX_194}"
    , 405 => "{INITX_195}"
    , 406 => "{INITX_196}"
    , 407 => "{INITX_197}"
    , 408 => "{INITX_198}"
    , 409 => "{INITX_199}"
    , 410 => "{INITX_19a}"
    , 411 => "{INITX_19b}"
    , 412 => "{INITX_19c}"
    , 413 => "{INITX_19d}"
    , 414 => "{INITX_19e}"
    , 415 => "{INITX_19f}"
    , 416 => "{INITX_1a0}"
    , 417 => "{INITX_1a1}"
    , 418 => "{INITX_1a2}"
    , 419 => "{INITX_1a3}"
    , 420 => "{INITX_1a4}"
    , 421 => "{INITX_1a5}"
    , 422 => "{INITX_1a6}"
    , 423 => "{INITX_1a7}"
    , 424 => "{INITX_1a8}"
    , 425 => "{INITX_1a9}"
    , 426 => "{INITX_1aa}"
    , 427 => "{INITX_1ab}"
    , 428 => "{INITX_1ac}"
    , 429 => "{INITX_1ad}"
    , 430 => "{INITX_1ae}"
    , 431 => "{INITX_1af}"
    , 432 => "{INITX_1b0}"
    , 433 => "{INITX_1b1}"
    , 434 => "{INITX_1b2}"
    , 435 => "{INITX_1b3}"
    , 436 => "{INITX_1b4}"
    , 437 => "{INITX_1b5}"
    , 438 => "{INITX_1b6}"
    , 439 => "{INITX_1b7}"
    , 440 => "{INITX_1b8}"
    , 441 => "{INITX_1b9}"
    , 442 => "{INITX_1ba}"
    , 443 => "{INITX_1bb}"
    , 444 => "{INITX_1bc}"
    , 445 => "{INITX_1bd}"
    , 446 => "{INITX_1be}"
    , 447 => "{INITX_1bf}"
    , 448 => "{INITX_1c0}"
    , 449 => "{INITX_1c1}"
    , 450 => "{INITX_1c2}"
    , 451 => "{INITX_1c3}"
    , 452 => "{INITX_1c4}"
    , 453 => "{INITX_1c5}"
    , 454 => "{INITX_1c6}"
    , 455 => "{INITX_1c7}"
    , 456 => "{INITX_1c8}"
    , 457 => "{INITX_1c9}"
    , 458 => "{INITX_1ca}"
    , 459 => "{INITX_1cb}"
    , 460 => "{INITX_1cc}"
    , 461 => "{INITX_1cd}"
    , 462 => "{INITX_1ce}"
    , 463 => "{INITX_1cf}"
    , 464 => "{INITX_1d0}"
    , 465 => "{INITX_1d1}"
    , 466 => "{INITX_1d2}"
    , 467 => "{INITX_1d3}"
    , 468 => "{INITX_1d4}"
    , 469 => "{INITX_1d5}"
    , 470 => "{INITX_1d6}"
    , 471 => "{INITX_1d7}"
    , 472 => "{INITX_1d8}"
    , 473 => "{INITX_1d9}"
    , 474 => "{INITX_1da}"
    , 475 => "{INITX_1db}"
    , 476 => "{INITX_1dc}"
    , 477 => "{INITX_1dd}"
    , 478 => "{INITX_1de}"
    , 479 => "{INITX_1df}"
    , 480 => "{INITX_1e0}"
    , 481 => "{INITX_1e1}"
    , 482 => "{INITX_1e2}"
    , 483 => "{INITX_1e3}"
    , 484 => "{INITX_1e4}"
    , 485 => "{INITX_1e5}"
    , 486 => "{INITX_1e6}"
    , 487 => "{INITX_1e7}"
    , 488 => "{INITX_1e8}"
    , 489 => "{INITX_1e9}"
    , 490 => "{INITX_1ea}"
    , 491 => "{INITX_1eb}"
    , 492 => "{INITX_1ec}"
    , 493 => "{INITX_1ed}"
    , 494 => "{INITX_1ee}"
    , 495 => "{INITX_1ef}"
    , 496 => "{INITX_1f0}"
    , 497 => "{INITX_1f1}"
    , 498 => "{INITX_1f2}"
    , 499 => "{INITX_1f3}"
    , 500 => "{INITX_1f4}"
    , 501 => "{INITX_1f5}"
    , 502 => "{INITX_1f6}"
    , 503 => "{INITX_1f7}"
    , 504 => "{INITX_1f8}"
    , 505 => "{INITX_1f9}"
    , 506 => "{INITX_1fa}"
    , 507 => "{INITX_1fb}"
    , 508 => "{INITX_1fc}"
    , 509 => "{INITX_1fd}"
    , 510 => "{INITX_1fe}"
    , 511 => "{INITX_1ff}"
    , 512 => "{INITX_200}"
    , 513 => "{INITX_201}"
    , 514 => "{INITX_202}"
    , 515 => "{INITX_203}"
    , 516 => "{INITX_204}"
    , 517 => "{INITX_205}"
    , 518 => "{INITX_206}"
    , 519 => "{INITX_207}"
    , 520 => "{INITX_208}"
    , 521 => "{INITX_209}"
    , 522 => "{INITX_20a}"
    , 523 => "{INITX_20b}"
    , 524 => "{INITX_20c}"
    , 525 => "{INITX_20d}"
    , 526 => "{INITX_20e}"
    , 527 => "{INITX_20f}"
    , 528 => "{INITX_210}"
    , 529 => "{INITX_211}"
    , 530 => "{INITX_212}"
    , 531 => "{INITX_213}"
    , 532 => "{INITX_214}"
    , 533 => "{INITX_215}"
    , 534 => "{INITX_216}"
    , 535 => "{INITX_217}"
    , 536 => "{INITX_218}"
    , 537 => "{INITX_219}"
    , 538 => "{INITX_21a}"
    , 539 => "{INITX_21b}"
    , 540 => "{INITX_21c}"
    , 541 => "{INITX_21d}"
    , 542 => "{INITX_21e}"
    , 543 => "{INITX_21f}"
    , 544 => "{INITX_220}"
    , 545 => "{INITX_221}"
    , 546 => "{INITX_222}"
    , 547 => "{INITX_223}"
    , 548 => "{INITX_224}"
    , 549 => "{INITX_225}"
    , 550 => "{INITX_226}"
    , 551 => "{INITX_227}"
    , 552 => "{INITX_228}"
    , 553 => "{INITX_229}"
    , 554 => "{INITX_22a}"
    , 555 => "{INITX_22b}"
    , 556 => "{INITX_22c}"
    , 557 => "{INITX_22d}"
    , 558 => "{INITX_22e}"
    , 559 => "{INITX_22f}"
    , 560 => "{INITX_230}"
    , 561 => "{INITX_231}"
    , 562 => "{INITX_232}"
    , 563 => "{INITX_233}"
    , 564 => "{INITX_234}"
    , 565 => "{INITX_235}"
    , 566 => "{INITX_236}"
    , 567 => "{INITX_237}"
    , 568 => "{INITX_238}"
    , 569 => "{INITX_239}"
    , 570 => "{INITX_23a}"
    , 571 => "{INITX_23b}"
    , 572 => "{INITX_23c}"
    , 573 => "{INITX_23d}"
    , 574 => "{INITX_23e}"
    , 575 => "{INITX_23f}"
    , 576 => "{INITX_240}"
    , 577 => "{INITX_241}"
    , 578 => "{INITX_242}"
    , 579 => "{INITX_243}"
    , 580 => "{INITX_244}"
    , 581 => "{INITX_245}"
    , 582 => "{INITX_246}"
    , 583 => "{INITX_247}"
    , 584 => "{INITX_248}"
    , 585 => "{INITX_249}"
    , 586 => "{INITX_24a}"
    , 587 => "{INITX_24b}"
    , 588 => "{INITX_24c}"
    , 589 => "{INITX_24d}"
    , 590 => "{INITX_24e}"
    , 591 => "{INITX_24f}"
    , 592 => "{INITX_250}"
    , 593 => "{INITX_251}"
    , 594 => "{INITX_252}"
    , 595 => "{INITX_253}"
    , 596 => "{INITX_254}"
    , 597 => "{INITX_255}"
    , 598 => "{INITX_256}"
    , 599 => "{INITX_257}"
    , 600 => "{INITX_258}"
    , 601 => "{INITX_259}"
    , 602 => "{INITX_25a}"
    , 603 => "{INITX_25b}"
    , 604 => "{INITX_25c}"
    , 605 => "{INITX_25d}"
    , 606 => "{INITX_25e}"
    , 607 => "{INITX_25f}"
    , 608 => "{INITX_260}"
    , 609 => "{INITX_261}"
    , 610 => "{INITX_262}"
    , 611 => "{INITX_263}"
    , 612 => "{INITX_264}"
    , 613 => "{INITX_265}"
    , 614 => "{INITX_266}"
    , 615 => "{INITX_267}"
    , 616 => "{INITX_268}"
    , 617 => "{INITX_269}"
    , 618 => "{INITX_26a}"
    , 619 => "{INITX_26b}"
    , 620 => "{INITX_26c}"
    , 621 => "{INITX_26d}"
    , 622 => "{INITX_26e}"
    , 623 => "{INITX_26f}"
    , 624 => "{INITX_270}"
    , 625 => "{INITX_271}"
    , 626 => "{INITX_272}"
    , 627 => "{INITX_273}"
    , 628 => "{INITX_274}"
    , 629 => "{INITX_275}"
    , 630 => "{INITX_276}"
    , 631 => "{INITX_277}"
    , 632 => "{INITX_278}"
    , 633 => "{INITX_279}"
    , 634 => "{INITX_27a}"
    , 635 => "{INITX_27b}"
    , 636 => "{INITX_27c}"
    , 637 => "{INITX_27d}"
    , 638 => "{INITX_27e}"
    , 639 => "{INITX_27f}"
    , 640 => "{INITX_280}"
    , 641 => "{INITX_281}"
    , 642 => "{INITX_282}"
    , 643 => "{INITX_283}"
    , 644 => "{INITX_284}"
    , 645 => "{INITX_285}"
    , 646 => "{INITX_286}"
    , 647 => "{INITX_287}"
    , 648 => "{INITX_288}"
    , 649 => "{INITX_289}"
    , 650 => "{INITX_28a}"
    , 651 => "{INITX_28b}"
    , 652 => "{INITX_28c}"
    , 653 => "{INITX_28d}"
    , 654 => "{INITX_28e}"
    , 655 => "{INITX_28f}"
    , 656 => "{INITX_290}"
    , 657 => "{INITX_291}"
    , 658 => "{INITX_292}"
    , 659 => "{INITX_293}"
    , 660 => "{INITX_294}"
    , 661 => "{INITX_295}"
    , 662 => "{INITX_296}"
    , 663 => "{INITX_297}"
    , 664 => "{INITX_298}"
    , 665 => "{INITX_299}"
    , 666 => "{INITX_29a}"
    , 667 => "{INITX_29b}"
    , 668 => "{INITX_29c}"
    , 669 => "{INITX_29d}"
    , 670 => "{INITX_29e}"
    , 671 => "{INITX_29f}"
    , 672 => "{INITX_2a0}"
    , 673 => "{INITX_2a1}"
    , 674 => "{INITX_2a2}"
    , 675 => "{INITX_2a3}"
    , 676 => "{INITX_2a4}"
    , 677 => "{INITX_2a5}"
    , 678 => "{INITX_2a6}"
    , 679 => "{INITX_2a7}"
    , 680 => "{INITX_2a8}"
    , 681 => "{INITX_2a9}"
    , 682 => "{INITX_2aa}"
    , 683 => "{INITX_2ab}"
    , 684 => "{INITX_2ac}"
    , 685 => "{INITX_2ad}"
    , 686 => "{INITX_2ae}"
    , 687 => "{INITX_2af}"
    , 688 => "{INITX_2b0}"
    , 689 => "{INITX_2b1}"
    , 690 => "{INITX_2b2}"
    , 691 => "{INITX_2b3}"
    , 692 => "{INITX_2b4}"
    , 693 => "{INITX_2b5}"
    , 694 => "{INITX_2b6}"
    , 695 => "{INITX_2b7}"
    , 696 => "{INITX_2b8}"
    , 697 => "{INITX_2b9}"
    , 698 => "{INITX_2ba}"
    , 699 => "{INITX_2bb}"
    , 700 => "{INITX_2bc}"
    , 701 => "{INITX_2bd}"
    , 702 => "{INITX_2be}"
    , 703 => "{INITX_2bf}"
    , 704 => "{INITX_2c0}"
    , 705 => "{INITX_2c1}"
    , 706 => "{INITX_2c2}"
    , 707 => "{INITX_2c3}"
    , 708 => "{INITX_2c4}"
    , 709 => "{INITX_2c5}"
    , 710 => "{INITX_2c6}"
    , 711 => "{INITX_2c7}"
    , 712 => "{INITX_2c8}"
    , 713 => "{INITX_2c9}"
    , 714 => "{INITX_2ca}"
    , 715 => "{INITX_2cb}"
    , 716 => "{INITX_2cc}"
    , 717 => "{INITX_2cd}"
    , 718 => "{INITX_2ce}"
    , 719 => "{INITX_2cf}"
    , 720 => "{INITX_2d0}"
    , 721 => "{INITX_2d1}"
    , 722 => "{INITX_2d2}"
    , 723 => "{INITX_2d3}"
    , 724 => "{INITX_2d4}"
    , 725 => "{INITX_2d5}"
    , 726 => "{INITX_2d6}"
    , 727 => "{INITX_2d7}"
    , 728 => "{INITX_2d8}"
    , 729 => "{INITX_2d9}"
    , 730 => "{INITX_2da}"
    , 731 => "{INITX_2db}"
    , 732 => "{INITX_2dc}"
    , 733 => "{INITX_2dd}"
    , 734 => "{INITX_2de}"
    , 735 => "{INITX_2df}"
    , 736 => "{INITX_2e0}"
    , 737 => "{INITX_2e1}"
    , 738 => "{INITX_2e2}"
    , 739 => "{INITX_2e3}"
    , 740 => "{INITX_2e4}"
    , 741 => "{INITX_2e5}"
    , 742 => "{INITX_2e6}"
    , 743 => "{INITX_2e7}"
    , 744 => "{INITX_2e8}"
    , 745 => "{INITX_2e9}"
    , 746 => "{INITX_2ea}"
    , 747 => "{INITX_2eb}"
    , 748 => "{INITX_2ec}"
    , 749 => "{INITX_2ed}"
    , 750 => "{INITX_2ee}"
    , 751 => "{INITX_2ef}"
    , 752 => "{INITX_2f0}"
    , 753 => "{INITX_2f1}"
    , 754 => "{INITX_2f2}"
    , 755 => "{INITX_2f3}"
    , 756 => "{INITX_2f4}"
    , 757 => "{INITX_2f5}"
    , 758 => "{INITX_2f6}"
    , 759 => "{INITX_2f7}"
    , 760 => "{INITX_2f8}"
    , 761 => "{INITX_2f9}"
    , 762 => "{INITX_2fa}"
    , 763 => "{INITX_2fb}"
    , 764 => "{INITX_2fc}"
    , 765 => "{INITX_2fd}"
    , 766 => "{INITX_2fe}"
    , 767 => "{INITX_2ff}"
    , 768 => "{INITX_300}"
    , 769 => "{INITX_301}"
    , 770 => "{INITX_302}"
    , 771 => "{INITX_303}"
    , 772 => "{INITX_304}"
    , 773 => "{INITX_305}"
    , 774 => "{INITX_306}"
    , 775 => "{INITX_307}"
    , 776 => "{INITX_308}"
    , 777 => "{INITX_309}"
    , 778 => "{INITX_30a}"
    , 779 => "{INITX_30b}"
    , 780 => "{INITX_30c}"
    , 781 => "{INITX_30d}"
    , 782 => "{INITX_30e}"
    , 783 => "{INITX_30f}"
    , 784 => "{INITX_310}"
    , 785 => "{INITX_311}"
    , 786 => "{INITX_312}"
    , 787 => "{INITX_313}"
    , 788 => "{INITX_314}"
    , 789 => "{INITX_315}"
    , 790 => "{INITX_316}"
    , 791 => "{INITX_317}"
    , 792 => "{INITX_318}"
    , 793 => "{INITX_319}"
    , 794 => "{INITX_31a}"
    , 795 => "{INITX_31b}"
    , 796 => "{INITX_31c}"
    , 797 => "{INITX_31d}"
    , 798 => "{INITX_31e}"
    , 799 => "{INITX_31f}"
    , 800 => "{INITX_320}"
    , 801 => "{INITX_321}"
    , 802 => "{INITX_322}"
    , 803 => "{INITX_323}"
    , 804 => "{INITX_324}"
    , 805 => "{INITX_325}"
    , 806 => "{INITX_326}"
    , 807 => "{INITX_327}"
    , 808 => "{INITX_328}"
    , 809 => "{INITX_329}"
    , 810 => "{INITX_32a}"
    , 811 => "{INITX_32b}"
    , 812 => "{INITX_32c}"
    , 813 => "{INITX_32d}"
    , 814 => "{INITX_32e}"
    , 815 => "{INITX_32f}"
    , 816 => "{INITX_330}"
    , 817 => "{INITX_331}"
    , 818 => "{INITX_332}"
    , 819 => "{INITX_333}"
    , 820 => "{INITX_334}"
    , 821 => "{INITX_335}"
    , 822 => "{INITX_336}"
    , 823 => "{INITX_337}"
    , 824 => "{INITX_338}"
    , 825 => "{INITX_339}"
    , 826 => "{INITX_33a}"
    , 827 => "{INITX_33b}"
    , 828 => "{INITX_33c}"
    , 829 => "{INITX_33d}"
    , 830 => "{INITX_33e}"
    , 831 => "{INITX_33f}"
    , 832 => "{INITX_340}"
    , 833 => "{INITX_341}"
    , 834 => "{INITX_342}"
    , 835 => "{INITX_343}"
    , 836 => "{INITX_344}"
    , 837 => "{INITX_345}"
    , 838 => "{INITX_346}"
    , 839 => "{INITX_347}"
    , 840 => "{INITX_348}"
    , 841 => "{INITX_349}"
    , 842 => "{INITX_34a}"
    , 843 => "{INITX_34b}"
    , 844 => "{INITX_34c}"
    , 845 => "{INITX_34d}"
    , 846 => "{INITX_34e}"
    , 847 => "{INITX_34f}"
    , 848 => "{INITX_350}"
    , 849 => "{INITX_351}"
    , 850 => "{INITX_352}"
    , 851 => "{INITX_353}"
    , 852 => "{INITX_354}"
    , 853 => "{INITX_355}"
    , 854 => "{INITX_356}"
    , 855 => "{INITX_357}"
    , 856 => "{INITX_358}"
    , 857 => "{INITX_359}"
    , 858 => "{INITX_35a}"
    , 859 => "{INITX_35b}"
    , 860 => "{INITX_35c}"
    , 861 => "{INITX_35d}"
    , 862 => "{INITX_35e}"
    , 863 => "{INITX_35f}"
    , 864 => "{INITX_360}"
    , 865 => "{INITX_361}"
    , 866 => "{INITX_362}"
    , 867 => "{INITX_363}"
    , 868 => "{INITX_364}"
    , 869 => "{INITX_365}"
    , 870 => "{INITX_366}"
    , 871 => "{INITX_367}"
    , 872 => "{INITX_368}"
    , 873 => "{INITX_369}"
    , 874 => "{INITX_36a}"
    , 875 => "{INITX_36b}"
    , 876 => "{INITX_36c}"
    , 877 => "{INITX_36d}"
    , 878 => "{INITX_36e}"
    , 879 => "{INITX_36f}"
    , 880 => "{INITX_370}"
    , 881 => "{INITX_371}"
    , 882 => "{INITX_372}"
    , 883 => "{INITX_373}"
    , 884 => "{INITX_374}"
    , 885 => "{INITX_375}"
    , 886 => "{INITX_376}"
    , 887 => "{INITX_377}"
    , 888 => "{INITX_378}"
    , 889 => "{INITX_379}"
    , 890 => "{INITX_37a}"
    , 891 => "{INITX_37b}"
    , 892 => "{INITX_37c}"
    , 893 => "{INITX_37d}"
    , 894 => "{INITX_37e}"
    , 895 => "{INITX_37f}"
    , 896 => "{INITX_380}"
    , 897 => "{INITX_381}"
    , 898 => "{INITX_382}"
    , 899 => "{INITX_383}"
    , 900 => "{INITX_384}"
    , 901 => "{INITX_385}"
    , 902 => "{INITX_386}"
    , 903 => "{INITX_387}"
    , 904 => "{INITX_388}"
    , 905 => "{INITX_389}"
    , 906 => "{INITX_38a}"
    , 907 => "{INITX_38b}"
    , 908 => "{INITX_38c}"
    , 909 => "{INITX_38d}"
    , 910 => "{INITX_38e}"
    , 911 => "{INITX_38f}"
    , 912 => "{INITX_390}"
    , 913 => "{INITX_391}"
    , 914 => "{INITX_392}"
    , 915 => "{INITX_393}"
    , 916 => "{INITX_394}"
    , 917 => "{INITX_395}"
    , 918 => "{INITX_396}"
    , 919 => "{INITX_397}"
    , 920 => "{INITX_398}"
    , 921 => "{INITX_399}"
    , 922 => "{INITX_39a}"
    , 923 => "{INITX_39b}"
    , 924 => "{INITX_39c}"
    , 925 => "{INITX_39d}"
    , 926 => "{INITX_39e}"
    , 927 => "{INITX_39f}"
    , 928 => "{INITX_3a0}"
    , 929 => "{INITX_3a1}"
    , 930 => "{INITX_3a2}"
    , 931 => "{INITX_3a3}"
    , 932 => "{INITX_3a4}"
    , 933 => "{INITX_3a5}"
    , 934 => "{INITX_3a6}"
    , 935 => "{INITX_3a7}"
    , 936 => "{INITX_3a8}"
    , 937 => "{INITX_3a9}"
    , 938 => "{INITX_3aa}"
    , 939 => "{INITX_3ab}"
    , 940 => "{INITX_3ac}"
    , 941 => "{INITX_3ad}"
    , 942 => "{INITX_3ae}"
    , 943 => "{INITX_3af}"
    , 944 => "{INITX_3b0}"
    , 945 => "{INITX_3b1}"
    , 946 => "{INITX_3b2}"
    , 947 => "{INITX_3b3}"
    , 948 => "{INITX_3b4}"
    , 949 => "{INITX_3b5}"
    , 950 => "{INITX_3b6}"
    , 951 => "{INITX_3b7}"
    , 952 => "{INITX_3b8}"
    , 953 => "{INITX_3b9}"
    , 954 => "{INITX_3ba}"
    , 955 => "{INITX_3bb}"
    , 956 => "{INITX_3bc}"
    , 957 => "{INITX_3bd}"
    , 958 => "{INITX_3be}"
    , 959 => "{INITX_3bf}"
    , 960 => "{INITX_3c0}"
    , 961 => "{INITX_3c1}"
    , 962 => "{INITX_3c2}"
    , 963 => "{INITX_3c3}"
    , 964 => "{INITX_3c4}"
    , 965 => "{INITX_3c5}"
    , 966 => "{INITX_3c6}"
    , 967 => "{INITX_3c7}"
    , 968 => "{INITX_3c8}"
    , 969 => "{INITX_3c9}"
    , 970 => "{INITX_3ca}"
    , 971 => "{INITX_3cb}"
    , 972 => "{INITX_3cc}"
    , 973 => "{INITX_3cd}"
    , 974 => "{INITX_3ce}"
    , 975 => "{INITX_3cf}"
    , 976 => "{INITX_3d0}"
    , 977 => "{INITX_3d1}"
    , 978 => "{INITX_3d2}"
    , 979 => "{INITX_3d3}"
    , 980 => "{INITX_3d4}"
    , 981 => "{INITX_3d5}"
    , 982 => "{INITX_3d6}"
    , 983 => "{INITX_3d7}"
    , 984 => "{INITX_3d8}"
    , 985 => "{INITX_3d9}"
    , 986 => "{INITX_3da}"
    , 987 => "{INITX_3db}"
    , 988 => "{INITX_3dc}"
    , 989 => "{INITX_3dd}"
    , 990 => "{INITX_3de}"
    , 991 => "{INITX_3df}"
    , 992 => "{INITX_3e0}"
    , 993 => "{INITX_3e1}"
    , 994 => "{INITX_3e2}"
    , 995 => "{INITX_3e3}"
    , 996 => "{INITX_3e4}"
    , 997 => "{INITX_3e5}"
    , 998 => "{INITX_3e6}"
    , 999 => "{INITX_3e7}"
    ,1000 => "{INITX_3e8}"
    ,1001 => "{INITX_3e9}"
    ,1002 => "{INITX_3ea}"
    ,1003 => "{INITX_3eb}"
    ,1004 => "{INITX_3ec}"
    ,1005 => "{INITX_3ed}"
    ,1006 => "{INITX_3ee}"
    ,1007 => "{INITX_3ef}"
    ,1008 => "{INITX_3f0}"
    ,1009 => "{INITX_3f1}"
    ,1010 => "{INITX_3f2}"
    ,1011 => "{INITX_3f3}"
    ,1012 => "{INITX_3f4}"
    ,1013 => "{INITX_3f5}"
    ,1014 => "{INITX_3f6}"
    ,1015 => "{INITX_3f7}"
    ,1016 => "{INITX_3f8}"
    ,1017 => "{INITX_3f9}"
    ,1018 => "{INITX_3fa}"
    ,1019 => "{INITX_3fb}"
    ,1020 => "{INITX_3fc}"
    ,1021 => "{INITX_3fd}"
    ,1022 => "{INITX_3fe}"
    ,1023 => "{INITX_3ff}"
    );
  
begin

  process (clk_i) is
  begin  -- process
    if rising_edge(clk_i)
    then
      if (cke_i = '1')
      then
        instruction_o <= rom(conv_integer(address_i));
      end if;
    end if;
  end process;
  
--
end rom;

--
------------------------------------------------------------------------------------
--
-- END OF FILE {name}.vhd
--
------------------------------------------------------------------------------------

